





//parameter WIDTH=8;
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//    FILE Name     :  d_flip_flop.sv                                                                             //
//                                                                                                                //
//    Description   :  D ff will trasfer the Data when Reset is low                                               //
//                                                                                                                //
//    Inputs        :  clk,reset,D                                                                                //
//                                                                                                                //
//    Outputs       :  Q                                                                                          //
//                                                                                                                //
//
//                                                                                                                //
//                                                                                                                //
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////










module d_ff (
    input clk_i,
    input reset_i,
    input data_i,
    output reg q_o
);

  always @(posedge clk_i) begin
    if (reset_i) begin
      q_o <= 0;
    end  //      else if (D==1 || D ==0)  Q <=  D ;
    else begin
      q_o <= data_i;
    end
  end


endmodule

